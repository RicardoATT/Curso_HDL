module Mux_IP_Catalog(
	input 	A, B, C,
	output 	F);

MyMux u0(A, B, C, F);
 
endmodule 