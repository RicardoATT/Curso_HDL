
module MinionsII (
	clk_clk,
	leds_out_export,
	reset_reset_n);	

	input		clk_clk;
	output	[7:0]	leds_out_export;
	input		reset_reset_n;
endmodule
